module JumpCntTB();
    reg [1:0] j_type, branch_t;






endmodule